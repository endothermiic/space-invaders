module shots(clk, reset, keyPressed, xin, bulletX, bulletY, colour, drawEn);
//xin comes from output of rocket.v - xout from rocket.v 

input clk, reset, keyPressed;
wire updatePosEn, bulletActive, waitEn, topReached, userIntakeEn;
wire collidedWithAlien = 1'b0; //remove once aliens modulr working
input [7:0] xin;
output [7:0] bulletX;
output [6:0] bulletY; 
output [2:0] colour;
output drawEn;


datapathshot d0 (.clk(clk), .reset(reset), .updatePosEn(updatePosEn), .waitEn(waitEn), .xin(xin), .bulletX(bulletX),
					.bulletY(bulletY), .topReached(topReached), .colour(colour), .bulletActive(bulletActive));
controlpathshot c0 (.clk(clk), .reset(reset), .keyPressed(keyPressed), .topReached(topReached), .collidedWithAlien(collidedWithAlien),
	.updatedBulletPosition(bulletActive), .userIntakeEn(userIntakeEn), .updatePosEn(updatePosEn), .waitEn(waitEn), .drawEn(drawEn));

endmodule

module datapathshot(clk, reset, updatePosEn, waitEn, xin, bulletX, bulletY, topReached, bulletActive, colour);
	input clk, reset, updatePosEn, waitEn;
	input [7:0] xin; 
	wire [7:0] xinorig = xin;
	output reg [7:0] bulletX; 
	output reg [6:0] bulletY; 
//	reg [7:0] xout; 
//	reg [6:0] yout; 
	output reg [2:0] colour;
	output reg topReached, bulletActive;
	
	always @(posedge clk)
	begin
		if (~reset) 
			begin
				bulletX <= 8'd0; 
				bulletY <= 7'd105;
				topReached <= 1'b0;
				colour <= 3'b000;
				bulletActive <= 1'b0;
				topReached <= 1'b0;
			end
		else if (updatePosEn)
			begin
				bulletActive <= 1'b1;
				if (bulletY > 0) 
					begin
						bulletY <= bulletY - 5; //if not at top, move 5 units up - clear and redraw
						bulletX <= xinorig;
						colour <= 3'b111;
					end
				else begin
					bulletY <= 7'd105;
					bulletX <= xinorig;
					topReached <= 1'b1;
				end
			end
		else if (waitEn) colour <= 3'b000;
	end

	
endmodule



module controlpathshot (clk, reset, keyPressed, topReached, collidedWithAlien, updatedBulletPosition, userIntakeEn, updatePosEn, waitEn, drawEn);

	input clk, reset, keyPressed, topReached, collidedWithAlien, updatedBulletPosition;
	output reg userIntakeEn, updatePosEn, waitEn, drawEn;
	
	reg [2:0] current_state, next_state;
	
	localparam INTAKE = 2'd0, // Set frame counter for top boundary check to 0
				  //if bullet exists - erase it (ex if we reached top of screen or killed an alien)
												
					
				  UPDATE_POSITION = 2'd1, //update bullet position, draw bullet position, 
						          //pass the coordinates to the alienTalentManager back to check for collision
				  
				  WAIT = 2'd2; //check for collision, check for top reached, 
	

always @(*)
	begin: state_table
	
	case(current_state)
			INTAKE: next_state = (keyPressed) ? UPDATE_POSITION : INTAKE;
			
			UPDATE_POSITION: next_state = (collidedWithAlien || topReached) ? INTAKE : WAIT;
			
			WAIT: next_state = (updatedBulletPosition) ? UPDATE_POSITION : WAIT; 

		default: next_state = INTAKE;
	endcase
end

 
always @(*)
   begin: enable_signals
	
		userIntakeEn <= 1'b0;
		updatePosEn <= 1'b0;
		waitEn <= 1'b0;
	   drawEn <= 1'b0;
		
	case(current_state)
		INTAKE: userIntakeEn <= 1'b1;
		UPDATE_POSITION: begin updatePosEn <= 1'b1; drawEn <= 1'b1; end
		WAIT: waitEn <= 1'b1;
	endcase
		
end

//state transitions
always@(posedge clk)
	begin: state_transition
	if (~reset)
		begin
			current_state <= INTAKE;
		end
			
		else current_state <= next_state;
	end
endmodule
